-------------------------------------------------------------------------------
--
-- Title       : ALU
-- Design      : ProjectPartI
-- Author      : anirvan.kothuri@stonybrook.edu
-- Company     : Stony Brook University
--
-------------------------------------------------------------------------------
--
-- File        : C:
-- Generated   : Sun Oct 12 15:37:45 2025
-- From        : Interface description file
-- By          : ItfToHdl ver. 1.0
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--    and may be overwritten
--{entity {ALU} architecture {structural}}

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ALU is
	port(
		instr : in STD_LOGIC_VECTOR(5 downto 0);
		rs3 : out STD_LOGIC_VECTOR(127 downto 0)
		rs2 : out STD_LOGIC_VECTOR(127 downto 0)
		rs1 : out STD_LOGIC_VECTOR(127 downto 0)
		rd : out STD_LOGIC_VECTOR(127 downto 0);
	);
end ALU;

--}} End of automatically maintained section

architecture behavioral of ALU is
begin

	process(instr, rs3, rs2, rs1)
	begin
    	case instr
        	when "00000" =>    -- Load Immediate 
				case ld_in
			        when "000" => rd <= rd(127 downto 16) + imm;
			        when "001" => rd <= rd(127 downto 32) + imm + rd(15 downto 0);
			        when "010" => rd <= rd(127 downto 48) + imm + rd(31 downto 0);
			        when "011" => rd <= rd(127 downto 64) + imm + rd(47 downto 0);
			        when "100" => rd <= rd(127 downto 80) + imm + rd(63 downto 0);
			        when "101" => rd <= rd(127 downto 96) + imm + rd(79 downto 0);
			        when "110" => rd <= rd(127 downto 112) + imm + rd(95 downto 0);
			        when "111" => rd <= imm + rd(111 downto 0);

	        -- Multiply-Add and Multiply-Subtract R4-Instruction Format
	        when "00001" => -- Signed Integer Multiply-Add Low with Saturation 
	        when "00010" =>    -- Signed Integer Multiply-Add High with Saturation
	        when "00011" =>    -- Signed Integer Multiply-Subtract Low with Saturation
	        when "00100" =>    -- Signed Integer Multiply-Subtract High with Saturation
	        when "00101" =>    -- Signed Long Integer Multiply-Add Low with Saturation
	        when "00110" =>    -- Signed Long Integer Multiply-Add High with Saturation
	        when "00111" =>    -- Signed Long Integer Multiply-Subtract Low with Saturation
	        when "01000" =>    -- Signed Long Integer Multiply-Subtract High with Saturation
	
	        -- R3-Instruction Format
	        when "01001" =>    -- NOP
	        when "01010" =>    -- SHRHI
	        when "01011" =>    -- AU
	        when "01100" =>    -- CNT1H
	        when "01101" =>    -- AHS
	        when "01110" =>    -- OR
	        when "01111" =>    -- BCW
	        when "10000" =>    -- MAXWS
	        when "10001" =>    -- MINWS
	        when "10010" =>    -- MLHU
	        when "10011" =>    -- MLHCU
	        when "10100" =>    -- AND
	        when "10101" => -- CLZW
	        when "10110" =>    -- ROTW
	        when "10111" =>    -- SFWU
	        when "11000" =>    -- SFHS
		
			-- Invalid
			when others => 

end structural;	
